    others => (31 downto 0 => '0')
    );
end package rom;
